`define Q 8
`define PERIOD 20
